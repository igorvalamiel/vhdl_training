if operation = "0010" then
    c0 <= val1(0)*val2(0);
    c1 <= c0(val1(1)+val2(1)) + val1(1)*val2(1);
    c2 <= c0(val1(2)+val2(2)) + val1(2)*val2(2);
    c3 <= c0(val1(3)+val2(3)) + val1(3)*val2(3);
